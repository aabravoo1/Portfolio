module segment_15(in_x, ou_z);
	input [5:0] in_x;
	output reg[0:13] ou_z;
	
	parameter n0 = 6'b000000,
	          n1 = 6'b000001,
	          n2 = 6'b000010,
	          n3 = 6'b000011,
	          n4 = 6'b000100,
	          n5 = 6'b000101,
	          n6 = 6'b000110,
	          n7 = 6'b000111,
	          n8 = 6'b001000,
	          n9 = 6'b001001,
	          A  = 6'b001010,
	          B  = 6'b001011,
	          C  = 6'b001100,
	          D  = 6'b001101,
	          E  = 6'b001110,
	          F  = 6'b001111,
	          G  = 6'b010000,
	          H  = 6'b010001,
	          I  = 6'b010010,
	          J  = 6'b010011,
	          K  = 6'b010100,
	          L  = 6'b010101,
	          M  = 6'b010110,
	          N  = 6'b010111,
	          O  = 6'b011000,
	          P  = 6'b011001,
	          Q  = 6'b011010,
	          R  = 6'b011011,
	          S  = 6'b011100,
	          T  = 6'b011101,
	          U  = 6'b011110,
	          V  = 6'b011111,
	          W  = 6'b100000,
	          X  = 6'b100001,
	          Y  = 6'b100010,
	          Z  = 6'b100011;
	
	always @(in_x)
		begin
			case(in_x)
			n0 : ou_z = 14'b11111100000000;
			n1 : ou_z = 14'b01100000000000;
			n2 : ou_z = 14'b11011000011000;
			n3 : ou_z = 14'b11110000011000;
			n4 : ou_z = 14'b01100100011000;
			n5 : ou_z = 14'b10110100011000;
			n6 : ou_z = 14'b10111100011000;
			n7 : ou_z = 14'b11100000000000;
			n8 : ou_z = 14'b11111100011000;
			n9 : ou_z = 14'b11110100011000;
			A  : ou_z = 14'b11101100011000;
			B  : ou_z = 14'b11110001001010;
			C  : ou_z = 14'b10011100000000;
			D  : ou_z = 14'b11110001000010;
			E  : ou_z = 14'b10011100011000;
			F  : ou_z = 14'b10001100011000;
			G  : ou_z = 14'b10111100001111;
			H  : ou_z = 14'b01101100011000;
			I  : ou_z = 14'b10010001000010;
			J  : ou_z = 14'b01111000000000;
			K  : ou_z = 14'b00001100110001;
			L  : ou_z = 14'b00011100000000;
			M  : ou_z = 14'b01101110100000;
			N  : ou_z = 14'b01101110000001;
			O  : ou_z = 14'b11111100100100;
			P  : ou_z = 14'b11001100011000;
			Q  : ou_z = 14'b11111100000001;
			R  : ou_z = 14'b11001100011001;
			S  : ou_z = 14'b10110100011000;
			T  : ou_z = 14'b10000001000010;
			U  : ou_z = 14'b01111100000000;
			V  : ou_z = 14'b00001100100100;
			W  : ou_z = 14'b01101100000101;
			X  : ou_z = 14'b00000010100101;
			Y  : ou_z = 14'b01000100011010;
			Z  : ou_z = 14'b10010000100100;
	     default ou_z = 14'b00000000000000;
			endcase
		end
endmodule 
			
			
			
		
	
	