import mips_pkg::*;
module tb_multiplication;

localparam BIN_CODE_FILE="multiplication.txt";
localparam MULTIPLICAND = 5; // pos lim = 217   neg lim = 256 , -256
localparam MULTIPLIER   = -4; //pos lim = 151   neg lim = -128, 128
logic  clk;
logic  asyn_n_rst;

mips #(.FILE_NAME(BIN_CODE_FILE)) dut_mips(.*);

always begin
	clk = 0;
	#1ns;
	clk = 1;
	#1ns;
end

initial begin
	 tb_multiplication.dut_mips.dm_i.ram_mem[0] = MULTIPLICAND;
	 tb_multiplication.dut_mips.dm_i.ram_mem[1] = MULTIPLIER;
	 asyn_n_rst = 1;
	 #2ns;
	 asyn_n_rst = 0;
	 #2ns;
	 asyn_n_rst = 1; 
	 #2ns;

end

endmodule

/*
00010000000000010000000000000000
00010000000000100000000000000001
00101000000000110000000000000000
00010000000001000000000000000000
00001100010000100000000000000001
10001100010000000000000000001010
00000000100000010010000000100000
00001000011000110000000000000001
10000100010000110000000000000110
11000000000000000000000000010011
10001100001000000000000000001111
00000000100000010010000000100001
00001100011000110000000000000001
10000100010000110000000000001011
11000000000000000000000000010011
00001000010000100000000000000001
00000000100000010010000000100001
00001100011000110000000000000001
10000100010000110000000000010000
00010100000001000000000000000010
*/